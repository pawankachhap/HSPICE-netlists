Problem 3.52

D1 in out diode
C1 out 0 1u
R1 out 0 100
Vin in 0 SIN(0 5 60)

.model diode D
.tran 10n 100m
.end