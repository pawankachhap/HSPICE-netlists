High pass Filter example (AC response)
c1 in out 10p
r1 out 0 1k
vin in 0 ac 1
.ac dec 200 1meg 100meg
.end
